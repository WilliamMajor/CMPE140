
module compared(
    input wire [2:0] op,
    input wire [31:0] a, b,
    output wire zero
    );
    reg [31:0] y;
    assign zero = (y == 0);
    always @ (op, a, b) begin
        case (op)
            3'b000: y = a & b;
            3'b001: y = a | b;
            3'b010: y = a + b;
            3'b110: y = a - b;
            3'b111: y = (a < b) ? 1 : 0;
        endcase
    end
endmodule
